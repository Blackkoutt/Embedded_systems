module noise_generator (clk, enable, Q);
		input clk, enable;
		output [23:0] Q;
		reg [2:0] counter;
		
		always @(posedge clk)
			if (enable) counter = counter + 1'b1;
			
		assign Q = {{8{counter[2]}}, counter, 13'd0};
endmodule
