module product_generator(input [3:0] A, B,
								 output wire AB [3:0][3:0]);
					
	
	
endmodule
	
								 